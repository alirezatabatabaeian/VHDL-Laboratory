--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:07:25 10/03/2020
-- Design Name:   
-- Module Name:   E:/Proj/intro1/four1_test.vhd
-- Project Name:  intro1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: four_bit_adder
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY four1_test IS
END four1_test;
 
ARCHITECTURE behavior OF four1_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT four_bit_adder
    PORT(
         input1 : IN  std_logic_vector(3 downto 0);
         input2 : IN  std_logic_vector(3 downto 0);
         sub0 : IN  std_logic;
         output : OUT  std_logic_vector(4 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal input1 : std_logic_vector(3 downto 0) := (others => '0');
   signal input2 : std_logic_vector(3 downto 0) := (others => '0');
   signal sub0 : std_logic := '0';

 	--Outputs
   signal output : std_logic_vector(4 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
  
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: four_bit_adder PORT MAP (
          input1 => input1,
          input2 => input2,
          sub0 => sub0,
          output => output
        );

 

   -- Stimulus process
   stim_proc: process
   begin		
		sub0 <= '0';
		input1 <= "0000" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0000" ;
      input2 <= "1111" ;
		wait for 1 ns;

		input1 <= "0001" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0001" ;
      input2 <= "1111" ;
		wait for 1 ns;
 
		input1 <= "0010" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0010" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "0011" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0011" ;
      input2 <= "1111" ;
		wait for 1 ns;
      
		input1 <= "0100" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0100" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "0101" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0101" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "0110" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0110" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "0111" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "0111" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "1000" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1000" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "1001" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1001" ;
      input2 <= "1111" ;
		wait for 1 ns;
 
		input1 <= "1010" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1010" ;
      input2 <= "1111" ;
		wait for 1 ns;
	
		input1 <= "1011" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1011" ;
      input2 <= "1111" ;
		wait for 1 ns;
      
		input1 <= "1100" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1100" ;
      input2 <= "1111" ;
		wait for 1 ns;
	
		input1 <= "1101" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1101" ;
      input2 <= "1111" ;
		wait for 1 ns;
	
		input1 <= "1110" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1110" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
		input1 <= "1111" ;
      input2 <= "0000" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0001" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0011" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0100" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0101" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0110" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0111" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1000" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1001" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "0010" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1011" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1100" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1101" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1110" ;
		wait for 1 ns;
		input1 <= "1111" ;
      input2 <= "1111" ;
		wait for 1 ns;
		
      wait;
   end process;

END;
